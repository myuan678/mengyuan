class icache_down_transaction;
    import toy_pack::*;

    pc_req_t                            txreq;
    logic [MSHR_ENTRY_INDEX_WIDTH-1:0]  entry_id;
endclass:icache_down_transaction

