class icache_down_sequence;






endclass: icache_down_sequence
