// Lets say that the environment class was already there, and generator is
// a new component that needs to be included in the ENV.
class env;
  up_sequence 		        seq0; 			    // Generate transactions
  up_driver 			        d0; 			      // Driver to design
  up_monitor 			        m0; 			      // Monitor from design
  scoreboard 		          s0; 			      // Scoreboard connected to monitor
  mailbox 			          scb_mbx; 		    // Top level mailbox for SCB <-> MON
  virtual icache_up_if 	  icache_up_vif; 	// Virtual interface handle
  virtual icache_down_if 	icache_down_vif;

  event drv_done;
  mailbox drv_mbx;

  function new();
    d0 = new;
    m0 = new;
    s0 = new;
    scb_mbx = new();
    seq0 = new;
    drv_mbx = new;
  endfunction

  virtual task run();
    // Connect virtual interface handles
    d0.icache_up_vif = icache_up_vif;
    m0.icache_up_vif = icache_up_vif;
    d0.icache_down_vif = icache_down_vif;
    m0.icache_down_vif = icache_down_vif;

    // Connect mailboxes between each component
    d0.drv_mbx   = drv_mbx;
    seq0.drv_mbx = drv_mbx;

    m0.scb_mbx   = scb_mbx;
    s0.scb_mbx   = scb_mbx;

    // Connect event handles
    d0.drv_done   = drv_done;
    seq0.drv_done = drv_done;

    // Start all components - a fork join_any is used because
    // the stimulus is generated by the generator and we want the
    // simulation to exit only when the generator has finished
    // creating all transactions. Until then all other components
    // have to run in the background.
    fork
    	s0.run();
		d0.run();
    	m0.run();
      	seq0.run();
    join_any
  endtask
endclass