class icache_cfg;
    int pld_width = 32  ;
    bit debug_en  = 1   ;
endclass:icache_cfg